library verilog;
use verilog.vl_types.all;
entity Test_simtb is
end Test_simtb;
